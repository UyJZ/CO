`timescale 1ns / 1ps
module DREG(
    input clk,
	 input reset
    );


endmodule
